`ifdef word_width
`else
`define word_width 8
`endif

`ifdef stack_size
`else
`define stack_size 4
`endif
